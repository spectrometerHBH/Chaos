`timescale 1ns/1ps

`include "defines.v"

module PC(
    input wire clk, 
    input wire rst,


);
    
endmodule