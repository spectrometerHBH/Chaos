`timescale 1ns/1ps

`include "defines.v"

module PC(
    
);
    
endmodule